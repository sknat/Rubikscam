library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity VGA_OUT is
    port (
	 -- CLOCK
    CLOCK_25  : in std_logic;
	 -- material ports
    VGA_CLK   : out std_logic; --Clock
    VGA_HS    : out std_logic; --H_SYNC
    VGA_VS    : out std_logic; --V_SYNC
    VGA_BLANK : out std_logic; --BLANK
    VGA_SYNC  : out std_logic; --SYNC
    VGA_R     : out std_logic_vector(9 downto 0); --Red[9:0]
    VGA_G     : out std_logic_vector(9 downto 0); --Green[9:0]
    VGA_B     : out std_logic_vector(9 downto 0); --Blue[9:0]
	 -- program used ports
	 SCREEN_X  : out integer range 0 to 639 := 0;
	 SCREEN_Y  : out integer range 0 to 479 := 0;
	 VGA_DATA_R : in std_logic_vector(9 downto 0);
	 VGA_DATA_G : in std_logic_vector(9 downto 0);
	 VGA_DATA_B : in std_logic_vector(9 downto 0)
    );
end VGA_OUT;

architecture VGA_OUT_arch of VGA_OUT is

signal v_pos : integer range 0 to 524 := 0;
constant v_pixel_end : natural := 480;
constant v_sync_low : natural := 493;
constant v_sync_high : natural := 494;
constant v_end : natural := 524;


signal h_pos : integer range 0 to 799 := 0;
constant h_pixel_end : natural := 640;
constant h_sync_low : natural := 659;
constant h_sync_high : natural := 755;
constant h_end : natural := 799;


begin
process (CLOCK_25)
	begin
	 	if rising_edge(CLOCK_25) then
			--count pixels
			if h_pos < h_end then
				h_pos <= h_pos + 1;
			else
				-- end of line
				h_pos <= 0;
				if v_pos < v_end then
					v_pos <= v_pos + 1;
				else
					-- end of screen
					v_pos <= 0;
				end if;				
			end if;
			
			-- synchronisation signals generation
			if h_sync_low <= h_pos and h_pos <= h_sync_high then VGA_HS <= '0'; else VGA_HS <= '1'; end if;
			if v_sync_low <= v_pos and v_pos <= v_sync_high then VGA_VS <= '0'; else VGA_VS <= '1'; end if;
			
			-- update pixel
			if h_pos < h_pixel_end and v_pos < v_pixel_end then 
				VGA_B <= VGA_DATA_B;
				VGA_R <= VGA_DATA_R;
				VGA_G <= VGA_DATA_G;
				VGA_BLANK <= '1';
			else
				VGA_BLANK <= '0';
			end if;
			
		end if;
end process ;

SCREEN_X <= h_pos when h_pos < 640 else 0;
SCREEN_Y <= v_pos when v_pos < 480 else 0;

VGA_CLK <= CLOCK_25;
VGA_SYNC <= '0'; -- signal to keep to zero, overwise, synchronisation makes on green 

end VGA_OUT_arch;
